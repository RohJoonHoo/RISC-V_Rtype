`timescale 1ns / 1ps

module rom (
    input  logic [31:0] addr,
    output logic [31:0] data
);

logic [31:0]rom[0:15];

initial begin
    //rom[x] = 32'b func7_rs2_rs1_fnc3_rd_opcode; //R-Type
    rom[0] = 32'b0000000_00001_00010_000_00100_0110011; //add x4(23), x2(12), x1(11) 
    rom[1] = 32'b0100000_00001_00010_000_00101_0110011; //sub x5(1), x2(12), x1(11)
    rom[2] = 32'b0000000_00101_00010_001_00110_0110011; //SLL x6(24), x2(12), x5(1)
    rom[3] = 32'b0000000_00101_00010_101_00111_0110011; //SRL x7(6), x2(12), x5(1)
    rom[4] = 32'b0100000_00111_10000_101_01000_0110011; //SRA x8(ffc0_0000),x16(f000_0010),x7(d6)
    rom[5] = 32'b0000000_00001_10000_010_01001_0110011; //SLT x9(1),x16(f000_0010),x1('d11)
    rom[6] = 32'b0000000_10001_10000_010_01010_0110011; //SLT x10(1),x16(f000_0010),x17(f000_0011)
    rom[7] = 32'b0000000_00001_10000_011_01011_0110011; //SLTU x11(0),x16(f000_0010),x1('d11)
    rom[8] = 32'b0000000_00001_00010_100_01100_0110011; //XOR x12(7), x2(12), x1(11)
    rom[9] = 32'b0000000_00001_00010_110_01101_0110011; //OR x13(15), x2(12), x1(11)
    rom[10] = 32'b0000000_00001_00010_111_01110_0110011; //AND x14(8), x2(12), x1(11)
end

assign data = rom[addr[31:2]];

endmodule
